grammar edu:umn:cs:melt:exts:ableC:skeleton;

exports edu:umn:cs:melt:exts:ableC:skeleton:abstractsyntax;
exports edu:umn:cs:melt:exts:ableC:skeleton:concretesyntax;

